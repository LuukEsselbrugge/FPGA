-- barcodescanner_nios.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity barcodescanner_nios is
	port (
		clk_clk                             : in    std_logic                     := '0';             --                          clk.clk
		leds_external_connection_export     : out   std_logic_vector(7 downto 0);                     --     leds_external_connection.export
		ram_mem_odt                         : out   std_logic_vector(0 downto 0);                     --                          ram.mem_odt
		ram_mem_clk                         : inout std_logic_vector(0 downto 0)  := (others => '0'); --                             .mem_clk
		ram_mem_clk_n                       : inout std_logic_vector(0 downto 0)  := (others => '0'); --                             .mem_clk_n
		ram_mem_cs_n                        : out   std_logic_vector(0 downto 0);                     --                             .mem_cs_n
		ram_mem_cke                         : out   std_logic_vector(0 downto 0);                     --                             .mem_cke
		ram_mem_addr                        : out   std_logic_vector(12 downto 0);                    --                             .mem_addr
		ram_mem_ba                          : out   std_logic_vector(1 downto 0);                     --                             .mem_ba
		ram_mem_ras_n                       : out   std_logic;                                        --                             .mem_ras_n
		ram_mem_cas_n                       : out   std_logic;                                        --                             .mem_cas_n
		ram_mem_we_n                        : out   std_logic;                                        --                             .mem_we_n
		ram_mem_dq                          : inout std_logic_vector(7 downto 0)  := (others => '0'); --                             .mem_dq
		ram_mem_dqs                         : inout std_logic_vector(0 downto 0)  := (others => '0'); --                             .mem_dqs
		ram_mem_dm                          : out   std_logic_vector(0 downto 0);                     --                             .mem_dm
		ram_external_local_refresh_ack      : out   std_logic;                                        --                 ram_external.local_refresh_ack
		ram_external_local_init_done        : out   std_logic;                                        --                             .local_init_done
		ram_external_reset_phy_clk_n        : out   std_logic;                                        --                             .reset_phy_clk_n
		switches_external_connection_export : in    std_logic_vector(7 downto 0)  := (others => '0')  -- switches_external_connection.export
	);
end entity barcodescanner_nios;

architecture rtl of barcodescanner_nios is
	component barcodescanner_nios_ddr2_memory is
		port (
			local_address     : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			local_write_req   : in    std_logic                     := 'X';             -- write
			local_read_req    : in    std_logic                     := 'X';             -- read
			local_burstbegin  : in    std_logic                     := 'X';             -- beginbursttransfer
			local_ready       : out   std_logic;                                        -- waitrequest_n
			local_rdata       : out   std_logic_vector(15 downto 0);                    -- readdata
			local_rdata_valid : out   std_logic;                                        -- readdatavalid
			local_wdata       : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			local_be          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			local_size        : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			local_refresh_ack : out   std_logic;                                        -- export
			local_init_done   : out   std_logic;                                        -- export
			reset_phy_clk_n   : out   std_logic;                                        -- export
			mem_odt           : out   std_logic_vector(0 downto 0);                     -- mem_odt
			mem_clk           : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_clk
			mem_clk_n         : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_clk_n
			mem_cs_n          : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_cke           : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_addr          : out   std_logic_vector(12 downto 0);                    -- mem_addr
			mem_ba            : out   std_logic_vector(1 downto 0);                     -- mem_ba
			mem_ras_n         : out   std_logic;                                        -- mem_ras_n
			mem_cas_n         : out   std_logic;                                        -- mem_cas_n
			mem_we_n          : out   std_logic;                                        -- mem_we_n
			mem_dq            : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs           : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dm            : out   std_logic_vector(0 downto 0);                     -- mem_dm
			pll_ref_clk       : in    std_logic                     := 'X';             -- clk
			soft_reset_n      : in    std_logic                     := 'X';             -- reset_n
			global_reset_n    : in    std_logic                     := 'X';             -- reset_n
			reset_request_n   : out   std_logic;                                        -- reset_n
			phy_clk           : out   std_logic;                                        -- clk
			aux_full_rate_clk : out   std_logic;                                        -- clk
			aux_half_rate_clk : out   std_logic                                         -- clk
		);
	end component barcodescanner_nios_ddr2_memory;

	component barcodescanner_nios_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component barcodescanner_nios_jtag_uart_0;

	component barcodescanner_nios_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component barcodescanner_nios_leds;

	component barcodescanner_nios_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component barcodescanner_nios_nios2_gen2_0;

	component barcodescanner_nios_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component barcodescanner_nios_onchip_memory2_0;

	component barcodescanner_nios_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component barcodescanner_nios_switches;

	component barcodescanner_nios_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                               : in  std_logic                     := 'X';             -- clk
			ddr2_memory_sysclk_clk                                      : in  std_logic                     := 'X';             -- clk
			ddr2_memory_s1_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                        : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                               : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid                      : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                              : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                        : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                     : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid               : out std_logic;                                        -- readdatavalid
			ddr2_memory_s1_address                                      : out std_logic_vector(23 downto 0);                    -- address
			ddr2_memory_s1_write                                        : out std_logic;                                        -- write
			ddr2_memory_s1_read                                         : out std_logic;                                        -- read
			ddr2_memory_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			ddr2_memory_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			ddr2_memory_s1_beginbursttransfer                           : out std_logic;                                        -- beginbursttransfer
			ddr2_memory_s1_burstcount                                   : out std_logic_vector(2 downto 0);                     -- burstcount
			ddr2_memory_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			ddr2_memory_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			ddr2_memory_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                         : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                          : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    : out std_logic;                                        -- chipselect
			leds_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                               : out std_logic;                                        -- write
			leds_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                          : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                          : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                           : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                 : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                                   : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                   : out std_logic;                                        -- clken
			switches_s1_address                                         : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component barcodescanner_nios_mm_interconnect_0;

	component barcodescanner_nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component barcodescanner_nios_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_leds_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                              : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                 : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_switches_s1_readdata                          : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                   : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_ddr2_memory_s1_beginbursttransfer             : std_logic;                     -- mm_interconnect_0:ddr2_memory_s1_beginbursttransfer -> ddr2_memory:local_burstbegin
	signal mm_interconnect_0_ddr2_memory_s1_readdata                       : std_logic_vector(15 downto 0); -- ddr2_memory:local_rdata -> mm_interconnect_0:ddr2_memory_s1_readdata
	signal ddr2_memory_s1_waitrequest                                      : std_logic;                     -- ddr2_memory:local_ready -> ddr2_memory_s1_waitrequest:in
	signal mm_interconnect_0_ddr2_memory_s1_address                        : std_logic_vector(23 downto 0); -- mm_interconnect_0:ddr2_memory_s1_address -> ddr2_memory:local_address
	signal mm_interconnect_0_ddr2_memory_s1_read                           : std_logic;                     -- mm_interconnect_0:ddr2_memory_s1_read -> ddr2_memory:local_read_req
	signal mm_interconnect_0_ddr2_memory_s1_byteenable                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ddr2_memory_s1_byteenable -> ddr2_memory:local_be
	signal mm_interconnect_0_ddr2_memory_s1_readdatavalid                  : std_logic;                     -- ddr2_memory:local_rdata_valid -> mm_interconnect_0:ddr2_memory_s1_readdatavalid
	signal mm_interconnect_0_ddr2_memory_s1_write                          : std_logic;                     -- mm_interconnect_0:ddr2_memory_s1_write -> ddr2_memory:local_write_req
	signal mm_interconnect_0_ddr2_memory_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:ddr2_memory_s1_writedata -> ddr2_memory:local_wdata
	signal mm_interconnect_0_ddr2_memory_s1_burstcount                     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ddr2_memory_s1_burstcount -> ddr2_memory:local_size
	signal ddr2_memory_sysclk_clk                                          : std_logic;                     -- ddr2_memory:phy_clk -> mm_interconnect_0:ddr2_memory_sysclk_clk
	signal ddr2_memory_reset_request_n_reset                               : std_logic;                     -- ddr2_memory:reset_request_n -> ddr2_memory_reset_request_n_reset:in
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_ddr2_memory_s1_inv                            : std_logic;                     -- ddr2_memory_s1_waitrequest:inv -> mm_interconnect_0:ddr2_memory_s1_waitrequest
	signal ddr2_memory_reset_request_n_reset_ports_inv                     : std_logic;                     -- ddr2_memory_reset_request_n_reset:inv -> mm_interconnect_0:ddr2_memory_s1_translator_reset_reset_bridge_in_reset_reset
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [ddr2_memory:global_reset_n, ddr2_memory:soft_reset_n, jtag_uart_0:rst_n, leds:reset_n, nios2_gen2_0:reset_n, switches:reset_n]

begin

	ddr2_memory : component barcodescanner_nios_ddr2_memory
		port map (
			local_address     => mm_interconnect_0_ddr2_memory_s1_address,            --                  s1.address
			local_write_req   => mm_interconnect_0_ddr2_memory_s1_write,              --                    .write
			local_read_req    => mm_interconnect_0_ddr2_memory_s1_read,               --                    .read
			local_burstbegin  => mm_interconnect_0_ddr2_memory_s1_beginbursttransfer, --                    .beginbursttransfer
			local_ready       => ddr2_memory_s1_waitrequest,                          --                    .waitrequest_n
			local_rdata       => mm_interconnect_0_ddr2_memory_s1_readdata,           --                    .readdata
			local_rdata_valid => mm_interconnect_0_ddr2_memory_s1_readdatavalid,      --                    .readdatavalid
			local_wdata       => mm_interconnect_0_ddr2_memory_s1_writedata,          --                    .writedata
			local_be          => mm_interconnect_0_ddr2_memory_s1_byteenable,         --                    .byteenable
			local_size        => mm_interconnect_0_ddr2_memory_s1_burstcount,         --                    .burstcount
			local_refresh_ack => ram_external_local_refresh_ack,                      -- external_connection.export
			local_init_done   => ram_external_local_init_done,                        --                    .export
			reset_phy_clk_n   => ram_external_reset_phy_clk_n,                        --                    .export
			mem_odt           => ram_mem_odt,                                         --              memory.mem_odt
			mem_clk           => ram_mem_clk,                                         --                    .mem_clk
			mem_clk_n         => ram_mem_clk_n,                                       --                    .mem_clk_n
			mem_cs_n          => ram_mem_cs_n,                                        --                    .mem_cs_n
			mem_cke           => ram_mem_cke,                                         --                    .mem_cke
			mem_addr          => ram_mem_addr,                                        --                    .mem_addr
			mem_ba            => ram_mem_ba,                                          --                    .mem_ba
			mem_ras_n         => ram_mem_ras_n,                                       --                    .mem_ras_n
			mem_cas_n         => ram_mem_cas_n,                                       --                    .mem_cas_n
			mem_we_n          => ram_mem_we_n,                                        --                    .mem_we_n
			mem_dq            => ram_mem_dq,                                          --                    .mem_dq
			mem_dqs           => ram_mem_dqs,                                         --                    .mem_dqs
			mem_dm            => ram_mem_dm,                                          --                    .mem_dm
			pll_ref_clk       => clk_clk,                                             --              refclk.clk
			soft_reset_n      => rst_controller_reset_out_reset_ports_inv,            --        soft_reset_n.reset_n
			global_reset_n    => rst_controller_reset_out_reset_ports_inv,            --      global_reset_n.reset_n
			reset_request_n   => ddr2_memory_reset_request_n_reset,                   --     reset_request_n.reset_n
			phy_clk           => ddr2_memory_sysclk_clk,                              --              sysclk.clk
			aux_full_rate_clk => open,                                                --             auxfull.clk
			aux_half_rate_clk => open                                                 --             auxhalf.clk
		);

	jtag_uart_0 : component barcodescanner_nios_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	leds : component barcodescanner_nios_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	nios2_gen2_0 : component barcodescanner_nios_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component barcodescanner_nios_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	switches : component barcodescanner_nios_switches
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_external_connection_export       -- external_connection.export
		);

	mm_interconnect_0 : component barcodescanner_nios_mm_interconnect_0
		port map (
			clk_0_clk_clk                                               => clk_clk,                                                     --                                             clk_0_clk.clk
			ddr2_memory_sysclk_clk                                      => ddr2_memory_sysclk_clk,                                      --                                    ddr2_memory_sysclk.clk
			ddr2_memory_s1_translator_reset_reset_bridge_in_reset_reset => ddr2_memory_reset_request_n_reset_ports_inv,                 -- ddr2_memory_s1_translator_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                              --              nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                            => nios2_gen2_0_data_master_address,                            --                              nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                        => nios2_gen2_0_data_master_waitrequest,                        --                                                      .waitrequest
			nios2_gen2_0_data_master_byteenable                         => nios2_gen2_0_data_master_byteenable,                         --                                                      .byteenable
			nios2_gen2_0_data_master_read                               => nios2_gen2_0_data_master_read,                               --                                                      .read
			nios2_gen2_0_data_master_readdata                           => nios2_gen2_0_data_master_readdata,                           --                                                      .readdata
			nios2_gen2_0_data_master_readdatavalid                      => nios2_gen2_0_data_master_readdatavalid,                      --                                                      .readdatavalid
			nios2_gen2_0_data_master_write                              => nios2_gen2_0_data_master_write,                              --                                                      .write
			nios2_gen2_0_data_master_writedata                          => nios2_gen2_0_data_master_writedata,                          --                                                      .writedata
			nios2_gen2_0_data_master_debugaccess                        => nios2_gen2_0_data_master_debugaccess,                        --                                                      .debugaccess
			nios2_gen2_0_instruction_master_address                     => nios2_gen2_0_instruction_master_address,                     --                       nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                 => nios2_gen2_0_instruction_master_waitrequest,                 --                                                      .waitrequest
			nios2_gen2_0_instruction_master_read                        => nios2_gen2_0_instruction_master_read,                        --                                                      .read
			nios2_gen2_0_instruction_master_readdata                    => nios2_gen2_0_instruction_master_readdata,                    --                                                      .readdata
			nios2_gen2_0_instruction_master_readdatavalid               => nios2_gen2_0_instruction_master_readdatavalid,               --                                                      .readdatavalid
			ddr2_memory_s1_address                                      => mm_interconnect_0_ddr2_memory_s1_address,                    --                                        ddr2_memory_s1.address
			ddr2_memory_s1_write                                        => mm_interconnect_0_ddr2_memory_s1_write,                      --                                                      .write
			ddr2_memory_s1_read                                         => mm_interconnect_0_ddr2_memory_s1_read,                       --                                                      .read
			ddr2_memory_s1_readdata                                     => mm_interconnect_0_ddr2_memory_s1_readdata,                   --                                                      .readdata
			ddr2_memory_s1_writedata                                    => mm_interconnect_0_ddr2_memory_s1_writedata,                  --                                                      .writedata
			ddr2_memory_s1_beginbursttransfer                           => mm_interconnect_0_ddr2_memory_s1_beginbursttransfer,         --                                                      .beginbursttransfer
			ddr2_memory_s1_burstcount                                   => mm_interconnect_0_ddr2_memory_s1_burstcount,                 --                                                      .burstcount
			ddr2_memory_s1_byteenable                                   => mm_interconnect_0_ddr2_memory_s1_byteenable,                 --                                                      .byteenable
			ddr2_memory_s1_readdatavalid                                => mm_interconnect_0_ddr2_memory_s1_readdatavalid,              --                                                      .readdatavalid
			ddr2_memory_s1_waitrequest                                  => mm_interconnect_0_ddr2_memory_s1_inv,                        --                                                      .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --                         jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                                      .write
			jtag_uart_0_avalon_jtag_slave_read                          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                                      .read
			jtag_uart_0_avalon_jtag_slave_readdata                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                                      .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                                      .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                                      .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                                      .chipselect
			leds_s1_address                                             => mm_interconnect_0_leds_s1_address,                           --                                               leds_s1.address
			leds_s1_write                                               => mm_interconnect_0_leds_s1_write,                             --                                                      .write
			leds_s1_readdata                                            => mm_interconnect_0_leds_s1_readdata,                          --                                                      .readdata
			leds_s1_writedata                                           => mm_interconnect_0_leds_s1_writedata,                         --                                                      .writedata
			leds_s1_chipselect                                          => mm_interconnect_0_leds_s1_chipselect,                        --                                                      .chipselect
			nios2_gen2_0_debug_mem_slave_address                        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --                          nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                                      .write
			nios2_gen2_0_debug_mem_slave_read                           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                                      .read
			nios2_gen2_0_debug_mem_slave_readdata                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                                      .readdata
			nios2_gen2_0_debug_mem_slave_writedata                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                                      .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                                      .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                                      .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                                      .debugaccess
			onchip_memory2_0_s1_address                                 => mm_interconnect_0_onchip_memory2_0_s1_address,               --                                   onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                   => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                                      .write
			onchip_memory2_0_s1_readdata                                => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                                      .readdata
			onchip_memory2_0_s1_writedata                               => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                                      .writedata
			onchip_memory2_0_s1_byteenable                              => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                                      .byteenable
			onchip_memory2_0_s1_chipselect                              => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                                      .chipselect
			onchip_memory2_0_s1_clken                                   => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                                      .clken
			switches_s1_address                                         => mm_interconnect_0_switches_s1_address,                       --                                           switches_s1.address
			switches_s1_readdata                                        => mm_interconnect_0_switches_s1_readdata                       --                                                      .readdata
		);

	irq_mapper : component barcodescanner_nios_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_ddr2_memory_s1_inv <= not ddr2_memory_s1_waitrequest;

	ddr2_memory_reset_request_n_reset_ports_inv <= not ddr2_memory_reset_request_n_reset;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of barcodescanner_nios
