// barcodescanner_nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module barcodescanner_nios (
		input  wire        clk_clk,                                 //                                 clk.clk
		output wire        eth_tse_mac_mdio_connection_mdc,         //         eth_tse_mac_mdio_connection.mdc
		input  wire        eth_tse_mac_mdio_connection_mdio_in,     //                                    .mdio_in
		output wire        eth_tse_mac_mdio_connection_mdio_out,    //                                    .mdio_out
		output wire        eth_tse_mac_mdio_connection_mdio_oen,    //                                    .mdio_oen
		input  wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_in,   //        eth_tse_mac_rgmii_connection.rgmii_in
		output wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_out,  //                                    .rgmii_out
		input  wire        eth_tse_mac_rgmii_connection_rx_control, //                                    .rx_control
		output wire        eth_tse_mac_rgmii_connection_tx_control, //                                    .tx_control
		input  wire        eth_tse_mac_status_connection_set_10,    //       eth_tse_mac_status_connection.set_10
		input  wire        eth_tse_mac_status_connection_set_1000,  //                                    .set_1000
		output wire        eth_tse_mac_status_connection_eth_mode,  //                                    .eth_mode
		output wire        eth_tse_mac_status_connection_ena_10,    //                                    .ena_10
		input  wire        eth_tse_pcs_mac_rx_clock_connection_clk, // eth_tse_pcs_mac_rx_clock_connection.clk
		input  wire        eth_tse_pcs_mac_tx_clock_connection_clk, // eth_tse_pcs_mac_tx_clock_connection.clk
		input  wire [7:0]  pixelb_export,                           //                              pixelb.export
		input  wire [7:0]  pixelg_export,                           //                              pixelg.export
		input  wire [7:0]  pixelr_export,                           //                              pixelr.export
		output wire [7:0]  pixelselect_export,                      //                         pixelselect.export
		input  wire        reset_reset_n,                           //                               reset.reset_n
		input  wire [7:0]  switches_export,                         //                            switches.export
		input  wire [11:0] videoram_address,                        //                            videoram.address
		input  wire        videoram_chipselect,                     //                                    .chipselect
		input  wire        videoram_clken,                          //                                    .clken
		input  wire        videoram_write,                          //                                    .write
		output wire [31:0] videoram_readdata,                       //                                    .readdata
		input  wire [31:0] videoram_writedata,                      //                                    .writedata
		input  wire [3:0]  videoram_byteenable                      //                                    .byteenable
	);

	wire         sgdma_tx_out_valid;                                        // sgdma_tx:out_valid -> eth_tse:ff_tx_wren
	wire  [31:0] sgdma_tx_out_data;                                         // sgdma_tx:out_data -> eth_tse:ff_tx_data
	wire         sgdma_tx_out_ready;                                        // eth_tse:ff_tx_rdy -> sgdma_tx:out_ready
	wire         sgdma_tx_out_startofpacket;                                // sgdma_tx:out_startofpacket -> eth_tse:ff_tx_sop
	wire         sgdma_tx_out_endofpacket;                                  // sgdma_tx:out_endofpacket -> eth_tse:ff_tx_eop
	wire         sgdma_tx_out_error;                                        // sgdma_tx:out_error -> eth_tse:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                        // sgdma_tx:out_empty -> eth_tse:ff_tx_mod
	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                             // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [20:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                         // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_waitrequest;                      // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                          // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                             // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire         sgdma_tx_descriptor_read_readdatavalid;                    // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                         // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_waitrequest;                      // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                          // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                             // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire         sgdma_rx_descriptor_read_readdatavalid;                    // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire         sgdma_tx_descriptor_write_waitrequest;                     // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_address;                         // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                           // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                       // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire         sgdma_rx_descriptor_write_waitrequest;                     // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_address;                         // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                           // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                       // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [20:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] sgdma_tx_m_read_readdata;                                  // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_waitrequest;                               // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                   // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                      // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire         sgdma_tx_m_read_readdatavalid;                             // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire         sgdma_rx_m_write_waitrequest;                              // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_address;                                  // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire   [3:0] sgdma_rx_m_write_byteenable;                               // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         sgdma_rx_m_write_write;                                    // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire  [31:0] sgdma_rx_m_write_writedata;                                // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_eth_tse_control_port_readdata;           // eth_tse:reg_data_out -> mm_interconnect_0:eth_tse_control_port_readdata
	wire         mm_interconnect_0_eth_tse_control_port_waitrequest;        // eth_tse:reg_busy -> mm_interconnect_0:eth_tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_eth_tse_control_port_address;            // mm_interconnect_0:eth_tse_control_port_address -> eth_tse:reg_addr
	wire         mm_interconnect_0_eth_tse_control_port_read;               // mm_interconnect_0:eth_tse_control_port_read -> eth_tse:reg_rd
	wire         mm_interconnect_0_eth_tse_control_port_write;              // mm_interconnect_0:eth_tse_control_port_write -> eth_tse:reg_wr
	wire  [31:0] mm_interconnect_0_eth_tse_control_port_writedata;          // mm_interconnect_0:eth_tse_control_port_writedata -> eth_tse:reg_data_in
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                 // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                   // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                    // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_read;                       // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire         mm_interconnect_0_sgdma_rx_csr_write;                      // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                  // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                 // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                   // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                    // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_read;                       // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire         mm_interconnect_0_sgdma_tx_csr_write;                      // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                  // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;          // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;       // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;           // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;              // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;             // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [16:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;         // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;           // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s1_address;            // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;         // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;              // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;          // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;              // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_0_videoram_s1_chipselect;                  // mm_interconnect_0:VideoRAM_s1_chipselect -> VideoRAM:chipselect
	wire  [31:0] mm_interconnect_0_videoram_s1_readdata;                    // VideoRAM:readdata -> mm_interconnect_0:VideoRAM_s1_readdata
	wire  [11:0] mm_interconnect_0_videoram_s1_address;                     // mm_interconnect_0:VideoRAM_s1_address -> VideoRAM:address
	wire   [3:0] mm_interconnect_0_videoram_s1_byteenable;                  // mm_interconnect_0:VideoRAM_s1_byteenable -> VideoRAM:byteenable
	wire         mm_interconnect_0_videoram_s1_write;                       // mm_interconnect_0:VideoRAM_s1_write -> VideoRAM:write
	wire  [31:0] mm_interconnect_0_videoram_s1_writedata;                   // mm_interconnect_0:VideoRAM_s1_writedata -> VideoRAM:writedata
	wire         mm_interconnect_0_videoram_s1_clken;                       // mm_interconnect_0:VideoRAM_s1_clken -> VideoRAM:clken
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                       // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                        // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire  [31:0] mm_interconnect_0_pio_1_s1_readdata;                       // pio_1:readdata -> mm_interconnect_0:pio_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_1_s1_address;                        // mm_interconnect_0:pio_1_s1_address -> pio_1:address
	wire         mm_interconnect_0_pio_2_s1_chipselect;                     // mm_interconnect_0:pio_2_s1_chipselect -> pio_2:chipselect
	wire  [31:0] mm_interconnect_0_pio_2_s1_readdata;                       // pio_2:readdata -> mm_interconnect_0:pio_2_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_2_s1_address;                        // mm_interconnect_0:pio_2_s1_address -> pio_2:address
	wire         mm_interconnect_0_pio_2_s1_write;                          // mm_interconnect_0:pio_2_s1_write -> pio_2:write_n
	wire  [31:0] mm_interconnect_0_pio_2_s1_writedata;                      // mm_interconnect_0:pio_2_s1_writedata -> pio_2:writedata
	wire  [31:0] mm_interconnect_0_pio_3_s1_readdata;                       // pio_3:readdata -> mm_interconnect_0:pio_3_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_3_s1_address;                        // mm_interconnect_0:pio_3_s1_address -> pio_3:address
	wire  [31:0] mm_interconnect_0_pio_4_s1_readdata;                       // pio_4:readdata -> mm_interconnect_0:pio_4_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_4_s1_address;                        // mm_interconnect_0:pio_4_s1_address -> pio_4:address
	wire         irq_mapper_receiver0_irq;                                  // sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_irq_irq;                                             // irq_mapper:sender_irq -> nios2:irq
	wire         eth_tse_receive_valid;                                     // eth_tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] eth_tse_receive_data;                                      // eth_tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         eth_tse_receive_ready;                                     // avalon_st_adapter:in_0_ready -> eth_tse:ff_rx_rdy
	wire         eth_tse_receive_startofpacket;                             // eth_tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         eth_tse_receive_endofpacket;                               // eth_tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] eth_tse_receive_error;                                     // eth_tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] eth_tse_receive_empty;                                     // eth_tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                             // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                              // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                             // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                     // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                       // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                             // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                             // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [VideoRAM:reset, avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, eth_tse:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, onchip_memory:reset, pio_0:reset_n, pio_1:reset_n, pio_2:reset_n, pio_3:reset_n, pio_4:reset_n, rst_translator:in_reset, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [VideoRAM:reset_req, descriptor_memory:reset_req, nios2:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                           // nios2:debug_reset_request -> rst_controller:reset_in1

	barcodescanner_nios_VideoRAM videoram (
		.address     (mm_interconnect_0_videoram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_videoram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_videoram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_videoram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_videoram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_videoram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_videoram_s1_byteenable), //       .byteenable
		.address2    (videoram_address),                         //     s2.address
		.chipselect2 (videoram_chipselect),                      //       .chipselect
		.clken2      (videoram_clken),                           //       .clken
		.write2      (videoram_write),                           //       .write
		.readdata2   (videoram_readdata),                        //       .readdata
		.writedata2  (videoram_writedata),                       //       .writedata
		.byteenable2 (videoram_byteenable),                      //       .byteenable
		.clk         (clk_clk),                                  //   clk1.clk
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	barcodescanner_nios_descriptor_memory descriptor_memory (
		.clk        (clk_clk),                                           //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	barcodescanner_nios_eth_tse eth_tse (
		.clk           (clk_clk),                                            // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                     //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_eth_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_eth_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_eth_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_eth_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_eth_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_eth_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (eth_tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (eth_tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (eth_tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (eth_tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (eth_tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (eth_tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (eth_tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                            //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                            //     transmit_clock_connection.clk
		.ff_rx_data    (eth_tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (eth_tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (eth_tse_receive_error),                              //                              .error
		.ff_rx_mod     (eth_tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (eth_tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (eth_tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (eth_tse_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                                  //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                           //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                                 //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                                 //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                                 //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                         //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                                 //                              .valid
		.mdc           (eth_tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (eth_tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (eth_tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (eth_tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.magic_wakeup  (),                                                   //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (),                                                   //                              .magic_sleep_n
		.ff_tx_crc_fwd (),                                                   //                              .ff_tx_crc_fwd
		.ff_tx_septy   (),                                                   //                              .ff_tx_septy
		.tx_ff_uflow   (),                                                   //                              .tx_ff_uflow
		.ff_tx_a_full  (),                                                   //                              .ff_tx_a_full
		.ff_tx_a_empty (),                                                   //                              .ff_tx_a_empty
		.rx_err_stat   (),                                                   //                              .rx_err_stat
		.rx_frm_type   (),                                                   //                              .rx_frm_type
		.ff_rx_dsav    (),                                                   //                              .ff_rx_dsav
		.ff_rx_a_full  (),                                                   //                              .ff_rx_a_full
		.ff_rx_a_empty ()                                                    //                              .ff_rx_a_empty
	);

	barcodescanner_nios_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	barcodescanner_nios_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	barcodescanner_nios_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	barcodescanner_nios_pio_0 pio_0 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_0_s1_readdata), //                    .readdata
		.in_port  (switches_export)                      // external_connection.export
	);

	barcodescanner_nios_pio_0 pio_1 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_1_s1_readdata), //                    .readdata
		.in_port  (pixelr_export)                        // external_connection.export
	);

	barcodescanner_nios_pio_2 pio_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_2_s1_readdata),   //                    .readdata
		.out_port   (pixelselect_export)                     // external_connection.export
	);

	barcodescanner_nios_pio_0 pio_3 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_3_s1_readdata), //                    .readdata
		.in_port  (pixelg_export)                        // external_connection.export
	);

	barcodescanner_nios_pio_0 pio_4 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_4_s1_readdata), //                    .readdata
		.in_port  (pixelb_export)                        // external_connection.export
	);

	barcodescanner_nios_sgdma_rx sgdma_rx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	barcodescanner_nios_sgdma_tx sgdma_tx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	barcodescanner_nios_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                         (clk_clk),                                                   //                       sys_clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address               (nios2_data_master_address),                                 //                 nios2_data_master.address
		.nios2_data_master_waitrequest           (nios2_data_master_waitrequest),                             //                                  .waitrequest
		.nios2_data_master_byteenable            (nios2_data_master_byteenable),                              //                                  .byteenable
		.nios2_data_master_read                  (nios2_data_master_read),                                    //                                  .read
		.nios2_data_master_readdata              (nios2_data_master_readdata),                                //                                  .readdata
		.nios2_data_master_write                 (nios2_data_master_write),                                   //                                  .write
		.nios2_data_master_writedata             (nios2_data_master_writedata),                               //                                  .writedata
		.nios2_data_master_debugaccess           (nios2_data_master_debugaccess),                             //                                  .debugaccess
		.nios2_instruction_master_address        (nios2_instruction_master_address),                          //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                      //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),                             //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),                         //                                  .readdata
		.sgdma_rx_descriptor_read_address        (sgdma_rx_descriptor_read_address),                          //          sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest    (sgdma_rx_descriptor_read_waitrequest),                      //                                  .waitrequest
		.sgdma_rx_descriptor_read_read           (sgdma_rx_descriptor_read_read),                             //                                  .read
		.sgdma_rx_descriptor_read_readdata       (sgdma_rx_descriptor_read_readdata),                         //                                  .readdata
		.sgdma_rx_descriptor_read_readdatavalid  (sgdma_rx_descriptor_read_readdatavalid),                    //                                  .readdatavalid
		.sgdma_rx_descriptor_write_address       (sgdma_rx_descriptor_write_address),                         //         sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest   (sgdma_rx_descriptor_write_waitrequest),                     //                                  .waitrequest
		.sgdma_rx_descriptor_write_write         (sgdma_rx_descriptor_write_write),                           //                                  .write
		.sgdma_rx_descriptor_write_writedata     (sgdma_rx_descriptor_write_writedata),                       //                                  .writedata
		.sgdma_rx_m_write_address                (sgdma_rx_m_write_address),                                  //                  sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest            (sgdma_rx_m_write_waitrequest),                              //                                  .waitrequest
		.sgdma_rx_m_write_byteenable             (sgdma_rx_m_write_byteenable),                               //                                  .byteenable
		.sgdma_rx_m_write_write                  (sgdma_rx_m_write_write),                                    //                                  .write
		.sgdma_rx_m_write_writedata              (sgdma_rx_m_write_writedata),                                //                                  .writedata
		.sgdma_tx_descriptor_read_address        (sgdma_tx_descriptor_read_address),                          //          sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest    (sgdma_tx_descriptor_read_waitrequest),                      //                                  .waitrequest
		.sgdma_tx_descriptor_read_read           (sgdma_tx_descriptor_read_read),                             //                                  .read
		.sgdma_tx_descriptor_read_readdata       (sgdma_tx_descriptor_read_readdata),                         //                                  .readdata
		.sgdma_tx_descriptor_read_readdatavalid  (sgdma_tx_descriptor_read_readdatavalid),                    //                                  .readdatavalid
		.sgdma_tx_descriptor_write_address       (sgdma_tx_descriptor_write_address),                         //         sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest   (sgdma_tx_descriptor_write_waitrequest),                     //                                  .waitrequest
		.sgdma_tx_descriptor_write_write         (sgdma_tx_descriptor_write_write),                           //                                  .write
		.sgdma_tx_descriptor_write_writedata     (sgdma_tx_descriptor_write_writedata),                       //                                  .writedata
		.sgdma_tx_m_read_address                 (sgdma_tx_m_read_address),                                   //                   sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest             (sgdma_tx_m_read_waitrequest),                               //                                  .waitrequest
		.sgdma_tx_m_read_read                    (sgdma_tx_m_read_read),                                      //                                  .read
		.sgdma_tx_m_read_readdata                (sgdma_tx_m_read_readdata),                                  //                                  .readdata
		.sgdma_tx_m_read_readdatavalid           (sgdma_tx_m_read_readdatavalid),                             //                                  .readdatavalid
		.descriptor_memory_s1_address            (mm_interconnect_0_descriptor_memory_s1_address),            //              descriptor_memory_s1.address
		.descriptor_memory_s1_write              (mm_interconnect_0_descriptor_memory_s1_write),              //                                  .write
		.descriptor_memory_s1_readdata           (mm_interconnect_0_descriptor_memory_s1_readdata),           //                                  .readdata
		.descriptor_memory_s1_writedata          (mm_interconnect_0_descriptor_memory_s1_writedata),          //                                  .writedata
		.descriptor_memory_s1_byteenable         (mm_interconnect_0_descriptor_memory_s1_byteenable),         //                                  .byteenable
		.descriptor_memory_s1_chipselect         (mm_interconnect_0_descriptor_memory_s1_chipselect),         //                                  .chipselect
		.descriptor_memory_s1_clken              (mm_interconnect_0_descriptor_memory_s1_clken),              //                                  .clken
		.eth_tse_control_port_address            (mm_interconnect_0_eth_tse_control_port_address),            //              eth_tse_control_port.address
		.eth_tse_control_port_write              (mm_interconnect_0_eth_tse_control_port_write),              //                                  .write
		.eth_tse_control_port_read               (mm_interconnect_0_eth_tse_control_port_read),               //                                  .read
		.eth_tse_control_port_readdata           (mm_interconnect_0_eth_tse_control_port_readdata),           //                                  .readdata
		.eth_tse_control_port_writedata          (mm_interconnect_0_eth_tse_control_port_writedata),          //                                  .writedata
		.eth_tse_control_port_waitrequest        (mm_interconnect_0_eth_tse_control_port_waitrequest),        //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.nios2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),           //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),             //                                  .write
		.nios2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),              //                                  .read
		.nios2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),          //                                  .readdata
		.nios2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),         //                                  .writedata
		.nios2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),        //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),       //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),       //                                  .debugaccess
		.onchip_memory_s1_address                (mm_interconnect_0_onchip_memory_s1_address),                //                  onchip_memory_s1.address
		.onchip_memory_s1_write                  (mm_interconnect_0_onchip_memory_s1_write),                  //                                  .write
		.onchip_memory_s1_readdata               (mm_interconnect_0_onchip_memory_s1_readdata),               //                                  .readdata
		.onchip_memory_s1_writedata              (mm_interconnect_0_onchip_memory_s1_writedata),              //                                  .writedata
		.onchip_memory_s1_byteenable             (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                  .byteenable
		.onchip_memory_s1_chipselect             (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                  .chipselect
		.onchip_memory_s1_clken                  (mm_interconnect_0_onchip_memory_s1_clken),                  //                                  .clken
		.pio_0_s1_address                        (mm_interconnect_0_pio_0_s1_address),                        //                          pio_0_s1.address
		.pio_0_s1_readdata                       (mm_interconnect_0_pio_0_s1_readdata),                       //                                  .readdata
		.pio_1_s1_address                        (mm_interconnect_0_pio_1_s1_address),                        //                          pio_1_s1.address
		.pio_1_s1_readdata                       (mm_interconnect_0_pio_1_s1_readdata),                       //                                  .readdata
		.pio_2_s1_address                        (mm_interconnect_0_pio_2_s1_address),                        //                          pio_2_s1.address
		.pio_2_s1_write                          (mm_interconnect_0_pio_2_s1_write),                          //                                  .write
		.pio_2_s1_readdata                       (mm_interconnect_0_pio_2_s1_readdata),                       //                                  .readdata
		.pio_2_s1_writedata                      (mm_interconnect_0_pio_2_s1_writedata),                      //                                  .writedata
		.pio_2_s1_chipselect                     (mm_interconnect_0_pio_2_s1_chipselect),                     //                                  .chipselect
		.pio_3_s1_address                        (mm_interconnect_0_pio_3_s1_address),                        //                          pio_3_s1.address
		.pio_3_s1_readdata                       (mm_interconnect_0_pio_3_s1_readdata),                       //                                  .readdata
		.pio_4_s1_address                        (mm_interconnect_0_pio_4_s1_address),                        //                          pio_4_s1.address
		.pio_4_s1_readdata                       (mm_interconnect_0_pio_4_s1_readdata),                       //                                  .readdata
		.sgdma_rx_csr_address                    (mm_interconnect_0_sgdma_rx_csr_address),                    //                      sgdma_rx_csr.address
		.sgdma_rx_csr_write                      (mm_interconnect_0_sgdma_rx_csr_write),                      //                                  .write
		.sgdma_rx_csr_read                       (mm_interconnect_0_sgdma_rx_csr_read),                       //                                  .read
		.sgdma_rx_csr_readdata                   (mm_interconnect_0_sgdma_rx_csr_readdata),                   //                                  .readdata
		.sgdma_rx_csr_writedata                  (mm_interconnect_0_sgdma_rx_csr_writedata),                  //                                  .writedata
		.sgdma_rx_csr_chipselect                 (mm_interconnect_0_sgdma_rx_csr_chipselect),                 //                                  .chipselect
		.sgdma_tx_csr_address                    (mm_interconnect_0_sgdma_tx_csr_address),                    //                      sgdma_tx_csr.address
		.sgdma_tx_csr_write                      (mm_interconnect_0_sgdma_tx_csr_write),                      //                                  .write
		.sgdma_tx_csr_read                       (mm_interconnect_0_sgdma_tx_csr_read),                       //                                  .read
		.sgdma_tx_csr_readdata                   (mm_interconnect_0_sgdma_tx_csr_readdata),                   //                                  .readdata
		.sgdma_tx_csr_writedata                  (mm_interconnect_0_sgdma_tx_csr_writedata),                  //                                  .writedata
		.sgdma_tx_csr_chipselect                 (mm_interconnect_0_sgdma_tx_csr_chipselect),                 //                                  .chipselect
		.VideoRAM_s1_address                     (mm_interconnect_0_videoram_s1_address),                     //                       VideoRAM_s1.address
		.VideoRAM_s1_write                       (mm_interconnect_0_videoram_s1_write),                       //                                  .write
		.VideoRAM_s1_readdata                    (mm_interconnect_0_videoram_s1_readdata),                    //                                  .readdata
		.VideoRAM_s1_writedata                   (mm_interconnect_0_videoram_s1_writedata),                   //                                  .writedata
		.VideoRAM_s1_byteenable                  (mm_interconnect_0_videoram_s1_byteenable),                  //                                  .byteenable
		.VideoRAM_s1_chipselect                  (mm_interconnect_0_videoram_s1_chipselect),                  //                                  .chipselect
		.VideoRAM_s1_clken                       (mm_interconnect_0_videoram_s1_clken)                        //                                  .clken
	);

	barcodescanner_nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	barcodescanner_nios_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (eth_tse_receive_data),                  //     in_0.data
		.in_0_valid          (eth_tse_receive_valid),                 //         .valid
		.in_0_ready          (eth_tse_receive_ready),                 //         .ready
		.in_0_startofpacket  (eth_tse_receive_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (eth_tse_receive_endofpacket),           //         .endofpacket
		.in_0_empty          (eth_tse_receive_empty),                 //         .empty
		.in_0_error          (eth_tse_receive_error),                 //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
